module add_test;

    // 定义输入和输出
    reg [31:0] A;
    reg [31:0] B;
    reg Cin;
    wire [31:0] Sum;
    wire Cout;

    // 创建32位加法器实例
    thirtytwo_bit_adder uut (
        .A(A),
        .B(B),
        .Cin(Cin),
        .Sum(Sum),
        .Cout(Cout)
    );

    // 初始化输入
    initial begin
        A = 32'b111111111111111111111111111111111; // 例如，A = 2^32 - 1
        B = 32'b111111111111111111111111111111111; // 例如，B = 2^32 - 1
        Cin = 1'b0;  // 例如，没有进位
        #10;        // 等待10个时钟周期

        // 更改输入
        A = 32'b000000000000000000000000000000000; // 例如，A = 0
        B = 32'b000000000000000000000000000000000; // 例如，B = 0
        Cin = 1'b0;  // 例如，没有进位
        #10;        // 等待10个时钟周期

        // 继续添加更多的测试案例...
